
`timescale 1 ns / 1 ps

    module MACC16
    (
        input clk,
        input rst,
        input [15:0] main,
        input [15:0] sub,
        input [31:0] scale,
        output [15:0] out
    );
        wire [47:0] pout;
        assign out = pout[31:16];

            // DSP48E2: 48-bit Multi-Functional Arithmetic Block
        // UltraScale
        // Xilinx HDL Language Template, version 2018.2
        DSP48E2 #(
            // Feature Control Attributes: Data Path Selection
            .AMULTSEL("A"), // Selects A input to multiplier (A, AD)
            .A_INPUT("DIRECT"), // Selects A input source, "DIRECT" (A port) or "CASCADE" (ACIN port)
            .BMULTSEL("B"), // Selects B input to multiplier (AD, B)
            .B_INPUT("DIRECT"), // Selects B input source, "DIRECT" (B port) or "CASCADE" (BCIN port)
            .PREADDINSEL("A"), // Selects input to pre-adder (A, B)
            .RND(48'h000000000000), // Rounding Constant
            .USE_MULT("MULTIPLY"), // Select multiplier usage (DYNAMIC, MULTIPLY, NONE)
            .USE_SIMD("ONE48"), // SIMD selection (FOUR12, ONE48, TWO24)
            .USE_WIDEXOR("FALSE"), // Use the Wide XOR function (FALSE, TRUE)
            .XORSIMD("XOR24_48_96"), // Mode of operation for the Wide XOR (XOR12, XOR24_48_96)
            // Pattern Detector Attributes: Pattern Detection Configuration
            .AUTORESET_PATDET("NO_RESET"), // NO_RESET, RESET_MATCH, RESET_NOT_MATCH
            .AUTORESET_PRIORITY("RESET"), // Priority of AUTORESET vs. CEP (CEP, RESET).
            .MASK(48'h3fffffffffff), // 48-bit mask value for pattern detect (1=ignore)
            .PATTERN(48'h000000000000), // 48-bit pattern match for pattern detect
            .SEL_MASK("MASK"), // C, MASK, ROUNDING_MODE1, ROUNDING_MODE2
            .SEL_PATTERN("PATTERN"), // Select pattern value (C, PATTERN)
            .USE_PATTERN_DETECT("NO_PATDET"), // Enable pattern detect (NO_PATDET, PATDET)
            // Programmable Inversion Attributes: Specifies built-in programmable inversion on specific pins
            .IS_ALUMODE_INVERTED(4'b0000), // Optional inversion for ALUMODE
            .IS_CARRYIN_INVERTED(1'b0), // Optional inversion for CARRYIN
            .IS_CLK_INVERTED(1'b0), // Optional inversion for CLK
            .IS_INMODE_INVERTED(5'b00000), // Optional inversion for INMODE
            .IS_OPMODE_INVERTED(9'b000000000), // Optional inversion for OPMODE
            .IS_RSTALLCARRYIN_INVERTED(1'b0), // Optional inversion for RSTALLCARRYIN
            .IS_RSTALUMODE_INVERTED(1'b0), // Optional inversion for RSTALUMODE
            .IS_RSTA_INVERTED(1'b0), // Optional inversion for RSTA
            .IS_RSTB_INVERTED(1'b0), // Optional inversion for RSTB
            .IS_RSTCTRL_INVERTED(1'b0), // Optional inversion for RSTCTRL
            .IS_RSTC_INVERTED(1'b0), // Optional inversion for RSTC
            .IS_RSTD_INVERTED(1'b0), // Optional inversion for RSTD
            .IS_RSTINMODE_INVERTED(1'b0), // Optional inversion for RSTINMODE
            .IS_RSTM_INVERTED(1'b0), // Optional inversion for RSTM
            .IS_RSTP_INVERTED(1'b0), // Optional inversion for RSTP
            // Register Control Attributes: Pipeline Register Configuration
            .ACASCREG(1), // Number of pipeline stages between A/ACIN and ACOUT (0-2)
            .ADREG(1), // Pipeline stages for pre-adder (0-1)
            .ALUMODEREG(1), // Pipeline stages for ALUMODE (0-1)
            .AREG(1), // Pipeline stages for A (0-2)
            .BCASCREG(1), // Number of pipeline stages between B/BCIN and BCOUT (0-2)
            .BREG(1), // Pipeline stages for B (0-2)
            .CARRYINREG(1), // Pipeline stages for CARRYIN (0-1)
            .CARRYINSELREG(1), // Pipeline stages for CARRYINSEL (0-1)
            .CREG(1), // Pipeline stages for C (0-1)
            .DREG(1), // Pipeline stages for D (0-1)
            .INMODEREG(1), // Pipeline stages for INMODE (0-1)
            .MREG(1), // Multiplier pipeline stages (0-1)
            .OPMODEREG(1), // Pipeline stages for OPMODE (0-1)
            .PREG(1) // Number of pipeline stages for P (0-1)
        )
        DSP48E2_inst (
            // Control outputs: Control Inputs/Status Bits
            //.OVERFLOW(OVERFLOW), // 1-bit output: Overflow in add/acc
            //.PATTERNBDETECT(PATTERNBDETECT), // 1-bit output: Pattern bar detect
            //.PATTERNDETECT(PATTERNDETECT), // 1-bit output: Pattern detect
            //.UNDERFLOW(UNDERFLOW), // 1-bit output: Underflow in add/acc
            // Data outputs: Data Ports
            .P(pout), // 48-bit output: Primary data
            // Control inputs: Control Inputs/Status Bits
            .ALUMODE(4'b0000), // 4-bit input: ALU control
            .CARRYINSEL(3'b000), // 3-bit input: Carry select
            .CLK(clk), // 1-bit input: Clock
            .INMODE(5'b00000), // 5-bit input: INMODE control
            .OPMODE(9'b11_000_01_01), // 9-bit input: Operation mode
            // Data inputs: Data Ports
            .A(scale[29:0]), // 30-bit input: A data
            .B({ {2{sub[15]}}, sub}), // 18-bit input: B data
            .C({ {16{main[15]}}, main, 16'b0 }), // 48-bit input: C data
            .CARRYIN(1'b0), // 1-bit input: Carry-in
            .D(28'b0), // 27-bit input: D data
            // Reset/Clock Enable inputs: Reset/Clock Enable Inputs
            .CEA1(1'b0), // 1-bit input: Clock enable for 1st stage AREG
            .CEA2(1'b1), // 1-bit input: Clock enable for 2nd stage AREG
            .CEAD(1'b1), // 1-bit input: Clock enable for ADREG
            .CEALUMODE(1'b1), // 1-bit input: Clock enable for ALUMODE
            .CEB1(1'b0), // 1-bit input: Clock enable for 1st stage BREG
            .CEB2(1'b1), // 1-bit input: Clock enable for 2nd stage BREG
            .CEC(1'b1), // 1-bit input: Clock enable for CREG
            .CECARRYIN(1'b1), // 1-bit input: Clock enable for CARRYINREG
            .CECTRL(1'b1), // 1-bit input: Clock enable for OPMODEREG and CARRYINSELREG
            .CED(1'b1), // 1-bit input: Clock enable for DREG
            .CEINMODE(1'b1), // 1-bit input: Clock enable for INMODEREG
            .CEM(1'b1), // 1-bit input: Clock enable for MREG
            .CEP(1'b1), // 1-bit input: Clock enable for PREG
            .RSTA(rst), // 1-bit input: Reset for AREG
            .RSTALLCARRYIN(rst), // 1-bit input: Reset for CARRYINREG
            .RSTALUMODE(rst), // 1-bit input: Reset for ALUMODEREG
            .RSTB(rst), // 1-bit input: Reset for BREG
            .RSTC(rst), // 1-bit input: Reset for CREG
            .RSTCTRL(rst), // 1-bit input: Reset for OPMODEREG and CARRYINSELREG
            .RSTD(rst), // 1-bit input: Reset for DREG and ADREG
            .RSTINMODE(rst), // 1-bit input: Reset for INMODEREG        
            .RSTM(rst), // 1-bit input: Reset for MREG
            .RSTP(rst) // 1-bit input: Reset for PREG
        );        

    endmodule


	module AXIReflection_v1_0 #
	(
		// Users to add parameters here
		parameter integer INITIAL_DELAY    = 12'd250,
        parameter integer INITIAL_SCALE    = 32'h0001_0000,
        parameter integer INITIAL_BYPASS   = 1'b0,
		
		parameter integer USE_URAM = 0,

		// User parameters ends
		// Do not modify the parameters beyond this line


		// Parameters of Axi Slave Bus Interface S00_AXI
		parameter integer C_S00_AXI_DATA_WIDTH	= 32,
		parameter integer C_S00_AXI_ADDR_WIDTH	= 4,

		// Parameters of Axi Slave Bus Interface RF_IN:RF_OUT
		parameter integer C_AXI_STREAM_TDATA_WIDTH	= 256
	)
	(
		// Users to add ports here
		// User ports ends
		// Do not modify the ports beyond this line

		// Ports of Axi Slave Bus Interface S00_AXI
		input wire  s00_axi_aclk,
		input wire  s00_axi_aresetn,
		input wire [C_S00_AXI_ADDR_WIDTH-1 : 0] s00_axi_awaddr,
		input wire [2 : 0] s00_axi_awprot,
		input wire  s00_axi_awvalid,
		output wire  s00_axi_awready,
		input wire [C_S00_AXI_DATA_WIDTH-1 : 0] s00_axi_wdata,
		input wire [(C_S00_AXI_DATA_WIDTH/8)-1 : 0] s00_axi_wstrb,
		input wire  s00_axi_wvalid,
		output wire  s00_axi_wready,
		output wire [1 : 0] s00_axi_bresp,
		output wire  s00_axi_bvalid,
		input wire  s00_axi_bready,
		input wire [C_S00_AXI_ADDR_WIDTH-1 : 0] s00_axi_araddr,
		input wire [2 : 0] s00_axi_arprot,
		input wire  s00_axi_arvalid,
		output wire  s00_axi_arready,
		output wire [C_S00_AXI_DATA_WIDTH-1 : 0] s00_axi_rdata,
		output wire [1 : 0] s00_axi_rresp,
		output wire  s00_axi_rvalid,
		input wire  s00_axi_rready,

		input wire  axis_aclk,
		input wire  axis_aresetn,

		// Ports of Axi Slave Bus Interface RF_IN
		output wire  rf_in_tready,
		input wire [C_AXI_STREAM_TDATA_WIDTH-1 : 0] rf_in_tdata,
		input wire  rf_in_tvalid,

		// Ports of Axi Master Bus Interface RF_OUT
		output wire  rf_out_tvalid,
		output wire [C_AXI_STREAM_TDATA_WIDTH-1 : 0] rf_out_tdata,
		input wire  rf_out_tready
	);
// Instantiation of Axi Bus Interface S00_AXI
	AXIReflection_v1_0_S00_AXI # ( 
	    .INITIAL_DELAY(INITIAL_DELAY),
	    .INITIAL_SCALE(INITIAL_SCALE),
	    .INITIAL_BYPASS(INITIAL_BYPASS),
		.C_S_AXI_DATA_WIDTH(C_S00_AXI_DATA_WIDTH),
		.C_S_AXI_ADDR_WIDTH(C_S00_AXI_ADDR_WIDTH)
	) AXIReflection_v1_0_S00_AXI_inst (
	    .delay(delay_axilite),
	    .scale(scale_axilite),
	    .bypass(bypass_axilite),
        .S_AXI_ACLK(s00_axi_aclk),
		.S_AXI_ARESETN(s00_axi_aresetn),
		.S_AXI_AWADDR(s00_axi_awaddr),
		.S_AXI_AWPROT(s00_axi_awprot),
		.S_AXI_AWVALID(s00_axi_awvalid),
		.S_AXI_AWREADY(s00_axi_awready),
		.S_AXI_WDATA(s00_axi_wdata),
		.S_AXI_WSTRB(s00_axi_wstrb),
		.S_AXI_WVALID(s00_axi_wvalid),
		.S_AXI_WREADY(s00_axi_wready),
		.S_AXI_BRESP(s00_axi_bresp),
		.S_AXI_BVALID(s00_axi_bvalid),
		.S_AXI_BREADY(s00_axi_bready),
		.S_AXI_ARADDR(s00_axi_araddr),
		.S_AXI_ARPROT(s00_axi_arprot),
		.S_AXI_ARVALID(s00_axi_arvalid),
		.S_AXI_ARREADY(s00_axi_arready),
		.S_AXI_RDATA(s00_axi_rdata),
		.S_AXI_RRESP(s00_axi_rresp),
		.S_AXI_RVALID(s00_axi_rvalid),
		.S_AXI_RREADY(s00_axi_rready)
	);

	// Add user logic here

    localparam N_URAM = C_AXI_STREAM_TDATA_WIDTH / 64;
    localparam N_BRAM = C_AXI_STREAM_TDATA_WIDTH / 64;
    localparam N_ADDR = USE_URAM ? 12 : 11;
    localparam N_DSP = C_AXI_STREAM_TDATA_WIDTH / 16;
    localparam MAX_ADDR = {N_ADDR{1'b1}};        

	// Add user logic here
	reg [N_ADDR-1:0] waddr;
	wire [N_ADDR-1:0] raddr;
	wire [7*N_URAM-1:0] unused;    
	wire axilite_valid;
    wire [31:0] delay_axilite;
    wire [31:0] delay_sync;
    reg [31:0] delay;
    wire [31:0] scale_axilite;
    wire [31:0] scale_sync;
    reg [31:0] scale;
    wire bypass_axilite;
    wire bypass_sync;
    reg bypass;
    reg delay_send;
    wire delay_recv;
	
	wire [C_AXI_STREAM_TDATA_WIDTH-1:0] din;
    wire [C_AXI_STREAM_TDATA_WIDTH-1 : 0] reflection;
    wire [C_AXI_STREAM_TDATA_WIDTH-1 : 0] out_data;
	
	reg [10:0] bringup_count;

    wire ready;
    wire [N_URAM - 1: 0] tvalid_out;
        
    wire [17:0] we;
    
    localparam WAIT = 3'd0;
    localparam INIT = 3'd1;
    localparam RUN = 3'd7;
    
    reg[2:0] state;
    
    reg[127:0] last_write;
    
	// Add user logic here
    xpm_cdc_handshake #(
        .DEST_EXT_HSK(0),
        .DEST_SYNC_FF(2),
        .INIT_SYNC_FF(0),
        .SIM_ASSERT_CHK(1),
        .SRC_SYNC_FF(2),
        .WIDTH(64))
        delay_handshake(
            .dest_clk(aclk),
            .dest_out({ delay_sync, scale_sync }),
            .dest_req(axilite_valid),
            .src_clk(s00_axi_aclk),
            .src_in({ delay_axilite, scale_axilite }),
            .src_send(delay_send),
            .src_rcv(delay_recv)
        );

    reg [31:0] last_delay_axilite;
    
    always @(posedge s00_axi_aclk)
    begin
        if (~s00_axi_aresetn) begin
            delay_send <= 1'b0;
            last_delay_axilite <= 32'b0;
        end else if (delay_send) begin
            delay_send <= ~delay_recv;
        end else if (~delay_recv && delay_axilite != last_delay_axilite) begin
            delay_send <= 1;
            last_delay_axilite <= delay_axilite;
        end
    end
    
    always @(posedge aclk) 
    begin
        if (axilite_valid) begin
            delay <= delay_sync;
            scale <= ~scale_sync + 1;
            bypass <= bypass_sync;
        end        
    end
    
    reg [2:0] tvalid;
    
    assign rf_in_tready = ready;
    
    assign ready = (state == RUN);
    assign din = (state == RUN) ? rf_in_tdata : {C_AXI_STREAM_TDATA_WIDTH{1'b0}};
    assign we = (state == INIT) ? 18'b0 : {18{1'b1}};

    assign raddr = waddr - delay;    

    always @(posedge axis_aclk)
    begin
        if (~axis_aresetn) begin
            bringup_count <= 100;
            state <= WAIT;
            waddr <= 0;
            tvalid <= 3'b0;
        end else
            case (state)
            WAIT: 
            begin
                if (bringup_count > 0) 
                    bringup_count <= bringup_count - 1;
                else
                    state <= INIT;        
            end 
            INIT:
            begin
                if (waddr == MAX_ADDR) begin
                    waddr <= delay;
                    state <= RUN;
                end else begin
                    waddr <= waddr + 1;
                end
            end
            RUN:
            begin
                tvalid <= { tvalid[1:0], &tvalid_out };
                waddr <= waddr + 1;
            end
            endcase    
    end
    
    genvar i;
    
    generate
        if (USE_URAM) 
        begin
            for (i = 0; i < N_URAM; i = i + 1)
            begin
                URAM288_BASE #(.AUTO_SLEEP_LATENCY(8),            // Latency requirement to enter sleep mode   
                          .AVG_CONS_INACTIVE_CYCLES(10),     // Average concecutive inactive cycles when is SLEEP mode for power
                                                             // estimation   
                          .BWE_MODE_A("PARITY_INDEPENDENT"), // Port A Byte write control   
                          .BWE_MODE_B("PARITY_INDEPENDENT"), // Port B Byte write control   
                          .EN_AUTO_SLEEP_MODE("FALSE"),      // Enable to automatically enter sleep mode   
                          .EN_ECC_RD_A("FALSE"),             // Port A ECC encoder   
                          .EN_ECC_RD_B("FALSE"),             // Port B ECC encoder   
                          .EN_ECC_WR_A("FALSE"),             // Port A ECC decoder   
                          .EN_ECC_WR_B("FALSE"),             // Port B ECC decoder   
                          .IREG_PRE_A("TRUE"),              // Optional Port A input pipeline registers   
                          .IREG_PRE_B("FALSE"),              // Optional Port B input pipeline registers   
                          .IS_CLK_INVERTED(1'b0),            // Optional inverter for CLK   
                          .IS_EN_A_INVERTED(1'b0),           // Optional inverter for Port A enable   
                          .IS_EN_B_INVERTED(1'b0),           // Optional inverter for Port B enable   
                          .IS_RDB_WR_A_INVERTED(1'b0),       // Optional inverter for Port A read/write select
                          .IS_RDB_WR_B_INVERTED(1'b0),       // Optional inverter for Port B read/write select   
                          .IS_RST_A_INVERTED(1'b0),          // Optional inverter for Port A reset   
                          .IS_RST_B_INVERTED(1'b0),          // Optional inverter for Port B reset   
                          .OREG_A("FALSE"),                  // Optional Port A output pipeline registers   
                          .OREG_B("TRUE"),                   // Optional Port B output pipeline registers   
                          .OREG_ECC_A("FALSE"),              // Port A ECC decoder output   
                          .OREG_ECC_B("FALSE"),              // Port B output ECC decoder   
                          //.REG_CAS_A("FALSE"),               // Optional Port A cascade register   
                          //.REG_CAS_B("FALSE"),               // Optional Port B cascade register   
                          .RST_MODE_A("ASYNC"),               // Port A reset mode   
                          .RST_MODE_B("ASYNC"),               // Port B reset mode   
                          //.SELF_ADDR_A(11'h000),             // Port A self-address value   
                          //.SELF_ADDR_B(11'h000),             // Port B self-address value   
                          //.SELF_MASK_A(11'h7ff),             // Port A self-address mask   
                          //.SELF_MASK_B(11'h7ff),             // Port B self-address mask   
                          .USE_EXT_CE_A("FALSE"),            // Enable Port A external CE inputs for output registers   
                          .USE_EXT_CE_B("FALSE")             // Enable Port B external CE inputs for output registers)
                    ) delay_data_fifo(.CLK(axis_aclk),
                    .ADDR_A({11'b0, waddr}), .ADDR_B({ 11'b0, raddr }), 
                    .BWE_A(we[8:0]), .BWE_B(9'h000),
                    .DIN_A({ 7'b0, rf_in_tvalid, din[64*i+:64] }), .DIN_B(71'h0),
                    /* .DOUT_A(), */ .DOUT_B({unused[7*i+:7], tvalid_out[i], reflection[64*i+:64]}),
                    .EN_A(state == RUN), .EN_B(state == RUN),
                    .INJECT_DBITERR_A(1'b0), .INJECT_DBITERR_B(1'b0),  
                    .INJECT_SBITERR_A(1'b0), .INJECT_SBITERR_B(1'b0),  
                    .OREG_CE_A(1'b0), .OREG_CE_B(1'b0),
                    .OREG_ECC_CE_A(1'b0),
                    .OREG_ECC_CE_B(1'b0),           // 1-bit input: Port B ECC decoder output register clock enable   
                    .RDB_WR_A(1'b1),                     // 1-bit input: Port A read/write select   
                    .RDB_WR_B(1'b0),                     // 1-bit input: Port B read/write select   
                    .RST_A(~axis_aresetn),            // 1-bit input: Port A asynchronous or synchronous reset for                                            
                                                             // output registers   
                    .RST_B(~axis_aresetn),           // 1-bit input: Port B asynchronous or synchronous reset for                                            
                                                             // output registers   
                    .SLEEP(1'b0)                            // 1-bit input: Dynamic power gating control
                    );
            end
        end else begin
            for (i = 0; i < N_BRAM; i = i + 1) 
            begin
                delay_fifo delay_data_fifo(.clka(axis_aclk),
                    .ena(state == RUN),
                    .wea(1'b1),
                    .addra(waddr),
                    .dina({rf_in_tvalid, din[64*i+:64]}),
                    .clkb(aclk),
                    .enb(state == RUN),
                    .addrb(raddr),
                    .doutb({tvalid_out[i], reflection[64*i+:64]}));
            end
        end

        for (i = 0; i < N_DSP; i = i + 1) begin
            MACC16 macc(.clk(axis_aclk), .rst(~axis_aresetn),
                .scale(scale),
                .main(ready ? rf_in_tdata[16*i+:16] : 16'b0), 
                .sub(ready ? reflection[16*i+:16] : 16'b0), 
                .out(out_data[16*i+:16]));
        end

    endgenerate        

    assign rf_out_tdata = bypass ? rf_in_tdata : out_data;
    assign rf_out_tvalid = ready & (bypass ? rf_in_tvalid : tvalid);
    

	// User logic ends

	endmodule
